`include "../mips_cpu.svh"

import mips_core_pkg::*;
